--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 


library IEEE;
use IEEE.STD_LOGIC_1164.all;

package pong_pack_2 is

	type tableau is array (2 downto 0) of std_logic_vector(8 downto 0);


end pong_pack_2;
